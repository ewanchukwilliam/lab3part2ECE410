------------------------------------------------------------------------
-- University  : University of Alberta
-- Course      : ECE 410
-- Project     : Lab 3
-- File        : data_memory.vhdl
-- Authors     : Antonio Alejandro Andara Lara
-- Date        : 23-Oct-2025
------------------------------------------------------------------------
-- Description  : 1 KB data memory with 32-bit read/write interface.
--                Supports synchronous writes and asynchronous reads.
------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY combined_mem IS
    PORT (
        clock      : IN STD_LOGIC;
        write_en   : IN STD_LOGIC;
        address    : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        write_data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        data       : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE rtl OF combined_mem IS

    -- Byte-addressable RAM
    TYPE memory_data IS ARRAY (0 TO 1023) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL RAM : memory_data := (
        -- Program (little-endian) - Simple test cases with 2 registers

        -- LOAD DATA: Load simple values from memory
        -- lw x1, 100(x0)    -- Load 16 into x1
        0 => x"83", 1 => x"20", 2 => x"40", 3 => x"06",
        -- lw x2, 104(x0)    -- Load -8 into x2
        4 => x"03", 5 => x"21", 6 => x"80", 7 => x"06",

        -- ARITHMETIC OPERATIONS
        -- add x3, x1, x2    -- x3 = 16 + (-8) = 8
        8 => x"B3", 9 => x"81", 10 => x"20", 11 => x"00",
        -- sub x4, x1, x2    -- x4 = 16 - (-8) = 24
        12 => x"33", 13 => x"82", 14 => x"20", 15 => x"40",

        -- IMMEDIATE OPERATIONS
        -- addi x5, x1, 4    -- x5 = 16 + 4 = 20
        16 => x"93", 17 => x"82", 18 => x"40", 19 => x"00",

        -- SHIFT OPERATIONS (using existing registers)
        -- srai x6, x1, 2    -- x6 = 16 >> 2 = 4 (positive shift)
        20 => x"13", 21 => x"D3", 22 => x"20", 23 => x"40",
        -- srai x7, x2, 1    -- x7 = -8 >> 1 = -4 (negative shift with sign extension)
        24 => x"93", 25 => x"53", 26 => x"11", 27 => x"40",

        -- STORE OPERATION
        -- sw x3, 108(x0)    -- Store x3 (8) to memory address 108
        28 => x"23", 29 => x"24", 30 => x"30", 31 => x"06",

        -- BRANCH NOT TAKEN
        -- beq x1, x2, 8     -- Compare 16 == -8? NO, don't branch
        32 => x"63", 33 => x"04", 34 => x"20", 35 => x"00",
        -- addi x8, x1, 1    -- x8 = 16 + 1 = 17 (this WILL execute)
        36 => x"13", 37 => x"04", 38 => x"11", 39 => x"00",

        -- BRANCH TAKEN
        -- beq x1, x1, 8     -- Compare 16 == 16? YES, branch
        40 => x"63", 41 => x"04", 42 => x"11", 43 => x"00",
        -- addi x9, x0, 99   -- x9 = 99 (this will be SKIPPED)
        44 => x"93", 45 => x"04", 46 => x"30", 47 => x"06",
        -- addi x9, x2, 2    -- x9 = -8 + 2 = -6 (this WILL execute after branch)
        48 => x"93", 49 => x"84", 50 => x"21", 51 => x"00",

        -- HALT
        52 => x"FF", 53 => x"FF", 54 => x"FF", 55 => x"FF",

        -- DATA SECTION
        100 => x"10", 101 => x"00", 102 => x"00", 103 => x"00",  -- 16
        104 => x"F8", 105 => x"FF", 106 => x"FF", 107 => x"FF",  -- -8 (0xFFFFFFF8)

        OTHERS => (OTHERS => '0')
    );

    SIGNAL addr_int : INTEGER := 0;

BEGIN
    addr_int <= to_integer(unsigned(address(9 DOWNTO 0))); -- Address conversion fits 1 KB

    PROCESS (clock)
    BEGIN
        IF rising_edge(clock) AND write_en = '1' THEN
            RAM(addr_int)     <= write_data(7 DOWNTO 0);
            RAM(addr_int + 1) <= write_data(15 DOWNTO 8);
            RAM(addr_int + 2) <= write_data(23 DOWNTO 16);
            RAM(addr_int + 3) <= write_data(31 DOWNTO 24);
        END IF;
    END PROCESS;

    -- read 4 consecutive bytes form one 32-bit word
    data <= RAM(addr_int + 3) &
        RAM(addr_int + 2) &
        RAM(addr_int + 1) &
        RAM(addr_int);

END ARCHITECTURE rtl;
